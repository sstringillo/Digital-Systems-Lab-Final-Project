module sprites(
	input logic clk,
	output logic [0:29][0:35][0:5] megaman_shooting_text,
	output logic [0:29][0:35][0:5] megaman_running1_text,
	output logic [0:29][0:35][0:5] megaman_running2_text,
	output logic [0:29][0:35][0:5] megaman_running3_text,
	output logic [0:29][0:35][0:5] megaman_jumping_text,
	output logic [0:27][0:26][0:5] soldier1_text,
	output logic [0:27][0:26][0:5] soldier2_text,
	output logic [0:28][0:34][0:5] soldierhigh1_text,
	output logic [0:28][0:34][0:5] soldierhigh2_text,
	output logic [0:34][0:88][0:5] tank1_text,
	output logic [0:34][0:88][0:5] tank2_text,
	output logic [0:34][0:88][0:5] tank3_text,
	output logic [0:29][0:35][0:5] boss_shooting_text,
	output logic [0:29][0:35][0:5] boss_running1_text,
	output logic [0:29][0:35][0:5] boss_running2_text,
	output logic [0:29][0:35][0:5] boss_running3_text,
	output logic [0:29][0:35][0:5] boss_jumping_text,
	output logic [0:2][0:5] bullet_text,
	output logic [0:1][0:2][0:5] rocket_text
);

always_comb
begin
//54 colors total, 6'hrepresented in 6 bits
megaman_shooting_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h10, 6'h10, 6'hf, 6'hf, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h15, 6'h1, 6'ha, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'h10, 6'hf, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'hf, 6'h1, 6'hf, 6'hf, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'h1, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h1, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'ha, 6'ha, 6'ha, 6'h1, 6'h15, 6'h34, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h34, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h34, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h11, 6'h11, 6'h11, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h1, 6'h12, 6'h12, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

megaman_running1_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h10, 6'h10, 6'hf, 6'hf, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'h10, 6'hf, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'ha, 6'ha, 6'h15, 6'h15, 6'h1, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'hf, 6'h1, 6'hf, 6'hf, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h1, 6'h1, 6'ha, 6'h11, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h1, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h1, 6'h15, 6'h15, 6'h34, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h12, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h34, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h12, 6'h12, 6'h12, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h12, 6'h12, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h12, 6'h12, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

megaman_running2_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h10, 6'h10, 6'hf, 6'hf, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'h10, 6'hf, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'hf, 6'h1, 6'hf, 6'hf, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'ha, 6'ha, 6'ha, 6'h1, 6'h11, 6'h11, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'h14, 6'h1, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h14, 6'h14, 6'h1, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h12, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

megaman_running3_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h10, 6'h10, 6'hf, 6'hf, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'h10, 6'hf, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'hf, 6'h1, 6'hf, 6'hf, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h11, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h11, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h15, 6'h1, 6'h1, 6'h1, 6'h15, 6'h1, 6'hf, 6'h1, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h12, 6'h14, 6'h14, 6'h14, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h12, 6'h12, 6'h12, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h12, 6'h12, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h1, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h12, 6'h12, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};
megaman_jumping_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h10, 6'h10, 6'hf, 6'hf, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h10, 6'h0},
'{6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'h15, 6'h1, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'hf, 6'h10, 6'hf, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'h2, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'hf, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'hf, 6'h1, 6'hf, 6'hf, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'h11, 6'h2, 6'h2, 6'h1, 6'h1, 6'ha, 6'h1, 6'h2, 6'ha, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h13, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'h11, 6'ha, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'hf, 6'h1, 6'h1, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h0, 6'hf, 6'hf, 6'hf, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h34, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h34, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h34, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h11, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h11, 6'h11, 6'h11, 6'h14, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h1, 6'h1, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h14, 6'h14, 6'h14, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};
soldier1_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h34, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h16, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h34, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2f, 6'h35, 6'h1, 6'h33, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h33, 6'h2f, 6'h1, 6'h2e, 6'h35, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h33, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h33, 6'h33, 6'h1, 6'h2e, 6'h35, 6'h35, 6'h2f, 6'h2f, 6'h35, 6'h35, 6'h35, 6'h33, 6'h33, 6'h1, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1d, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1, 6'h2f, 6'h2e, 6'h35, 6'h35, 6'h33, 6'h1d, 6'h1d, 6'h1d, 6'h2e, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h1f, 6'h1f, 6'h1, 6'h2f, 6'h2f, 6'h35, 6'h33, 6'h33, 6'h33, 6'h1, 6'h2e, 6'h2e, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h0, 6'h0, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2f, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h35, 6'h35, 6'h1, 6'h1, 6'h35, 6'h35, 6'h2f, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h35, 6'h1, 6'h33, 6'h33, 6'h1, 6'h35, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h35, 6'h1, 6'h33, 6'h2f, 6'h2f, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2f, 6'h2f, 6'h35, 6'h35, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h35, 6'h35, 6'h35, 6'h2e, 6'h33, 6'h33, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2e, 6'h2e, 6'h33, 6'h33, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h12, 6'h35, 6'h35, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0}
};
	
soldier2_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h34, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h16, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h34, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h1, 6'h1f, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2f, 6'h35, 6'h1, 6'h33, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h33, 6'h2f, 6'h1, 6'h2e, 6'h35, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h33, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h33, 6'h33, 6'h1, 6'h2e, 6'h35, 6'h35, 6'h2f, 6'h2f, 6'h35, 6'h35, 6'h35, 6'h33, 6'h33, 6'h1, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1d, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1d, 6'h1, 6'h2f, 6'h2e, 6'h35, 6'h35, 6'h33, 6'h1d, 6'h1d, 6'h1d, 6'h2e, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h1f, 6'h1f, 6'h1, 6'h2f, 6'h2f, 6'h35, 6'h33, 6'h33, 6'h33, 6'h1, 6'h2e, 6'h2e, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h0, 6'h0, 6'h1f, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2f, 6'h35, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h24, 6'h24, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h33, 6'h33, 6'h1, 6'h1, 6'h35, 6'h2e, 6'h2e, 6'h2f, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h33, 6'h1, 6'h2f, 6'h2f, 6'h1, 6'h35, 6'h33, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h35, 6'h1, 6'h2f, 6'h35, 6'h35, 6'h1, 6'h33, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h35, 6'h35, 6'h2f, 6'h2f, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2e, 6'h2e, 6'h1, 6'h2f, 6'h33, 6'h33, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2e, 6'h2e, 6'h35, 6'h1, 6'h2e, 6'h33, 6'h35, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h12, 6'h35, 6'h35, 6'h1, 6'h2e, 6'h35, 6'h35, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h12, 6'h12, 6'h12, 6'h12, 6'h1, 6'h12, 6'h12, 6'h12, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0}
};

soldierhigh1_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h1b, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h15, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1d, 6'h1d, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h15},
'{6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1f, 6'h1f, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1f, 6'h1d, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h0, 6'h15},
'{6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1f, 6'h1f, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h20, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h0, 6'h15},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h1, 6'h1, 6'h1f, 6'h1f, 6'h1, 6'h1e, 6'h20, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h15},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h1, 6'h1, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h19, 6'h1c, 6'h1a, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h1, 6'h20, 6'h20, 6'h1, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h19, 6'h19, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h19, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h19, 6'h19, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

soldierhigh2_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h21, 6'h1b, 6'h22, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'h1f, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h15, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1d, 6'h1d, 6'h1f, 6'h1f, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h15},
'{6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1f, 6'h1f, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h1, 6'h1f, 6'h1d, 6'h1d, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h0, 6'h15},
'{6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1f, 6'h1f, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h1, 6'h20, 6'h1, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1f, 6'h1, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h15, 6'h0, 6'h15},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h1, 6'h1, 6'h1f, 6'h1f, 6'h1, 6'h1e, 6'h20, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h15, 6'h15},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h1, 6'h1, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h19, 6'h1c, 6'h1a, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1e, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1e, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h1, 6'h20, 6'h20, 6'h1, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h20, 6'h20, 6'h20, 6'h20, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h20, 6'h20, 6'h1, 6'h20, 6'h20, 6'h20, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h19, 6'h19, 6'h19, 6'h1, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h19, 6'h19, 6'h19, 6'h1, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h19, 6'h19, 6'h19, 6'h19, 6'h1, 6'h19, 6'h19, 6'h19, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

tank1_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h1, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2c, 6'h1, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2d, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h28, 6'h1, 6'h25, 6'h25, 6'h29, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h28, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

tank2_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2c, 6'h1, 6'h2d, 6'h2d, 6'h2c, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h28, 6'h1, 6'h25, 6'h25, 6'h29, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h28, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

tank3_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h2c, 6'h1, 6'h2d, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h29, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2d, 6'h2d, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2d, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2d, 6'h2d, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h2c, 6'h29, 6'h29, 6'h0, 6'h0, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h26, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h1, 6'h1, 6'h1, 6'h25, 6'h25, 6'h25, 6'h25, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h24, 6'h28, 6'h1, 6'h25, 6'h25, 6'h29, 6'h29},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h25, 6'h25, 6'h25, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h29, 6'h29, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h29, 6'h25, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h2b, 6'h28, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h1, 6'h1, 6'h1, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h1, 6'h1, 6'h1, 6'h2b, 6'h28, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h29, 6'h1, 6'h28, 6'h28, 6'h28, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h2a, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h2b, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h1, 6'h26, 6'h27, 6'h27, 6'h2a, 6'h27, 6'h27, 6'h26, 6'h1, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h24, 6'h28, 6'h2b, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h27, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h28, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h27, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h26, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

boss_shooting_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'hc, 6'hb, 6'h2, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h3, 6'h3, 6'h5, 6'h5, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h3, 6'h5, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h3, 6'h3, 6'h8, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h3, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h9, 6'ha, 6'ha, 6'h9, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1}
};

boss_running1_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'hc, 6'hb, 6'h2, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h3, 6'h3, 6'h5, 6'h5, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'ha, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h3, 6'h5, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h3, 6'h3, 6'h8, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h3, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h9, 6'ha, 6'ha, 6'h9, 6'ha, 6'ha, 6'h1, 6'h1, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

boss_running2_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'hc, 6'hb, 6'h2, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h3, 6'h3, 6'h5, 6'h5, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'ha, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h3, 6'h5, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h3, 6'h3, 6'h8, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h3, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h9, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h1, 6'h4, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h1, 6'h4, 6'h4, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

boss_running3_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'hc, 6'hb, 6'h2, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h3, 6'h3, 6'h5, 6'h5, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h3, 6'h5, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h3, 6'h3, 6'h8, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h3, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h11, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h11, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

boss_jumping_text <=
'{
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0},
'{6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h5, 6'h3, 6'h3, 6'h5, 6'h5, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'hc, 6'hb, 6'h2, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h0, 6'h0, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0},
'{6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h3, 6'h5, 6'h3, 6'h0, 6'h0, 6'h0, 6'h1, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h6, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0},
'{6'h0, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h3, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'h2, 6'ha, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'h3, 6'h3, 6'h8, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h3, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'ha, 6'h2, 6'h7, 6'ha, 6'h7, 6'h7, 6'h2, 6'h2, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h2, 6'h2, 6'ha, 6'h2, 6'h2, 6'h2, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h8, 6'h8, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h1, 6'h1, 6'h1, 6'ha, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h9, 6'ha, 6'ha, 6'ha, 6'h9, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'ha, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'ha, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h4, 6'h4, 6'h4, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0},
'{6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h1, 6'h1, 6'h1, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0, 6'h0}
};

bullet_text <=
'{6'h17, 6'h17, 6'h17};

rocket_text <=
'{
'{6'h18, 6'h18, 6'h18},
'{6'h18, 6'h18, 6'h18}
};
end
endmodule

